library verilog;
use verilog.vl_types.all;
entity projectClock_vlg_vec_tst is
end projectClock_vlg_vec_tst;
